library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in  std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado     : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  	constant NOP  : std_logic_vector(3 downto 0) := "0000";
	constant LDA  : std_logic_vector(3 downto 0) := "0001";
	constant SOMA : std_logic_vector(3 downto 0) := "0010";
	constant SUB  : std_logic_vector(3 downto 0) := "0011";
	constant LDI  : std_logic_vector(3 downto 0) := "0100";
	constant STA  : std_logic_vector(3 downto 0) := "0101";
	constant JMP  : std_logic_vector(3 downto 0) := "0110";
	constant JSR  : std_logic_vector(3 downto 0) := "1001";
	constant RET  : std_logic_vector(3 downto 0) := "1010";
	constant JEQ  : std_logic_vector(3 downto 0) := "0111";
	constant CEQ  : std_logic_vector(3 downto 0) := "1000";

  
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

tmp(0) := NOP & '0' & x"00"; 	 ---- MAIN LOOP
tmp(1) := NOP & '0' & x"00"; 	 --%LABEL LOOP_INICIAL
tmp(2) := "1001000001110";	-- JSR @SR_INICIALIZACAO
tmp(3) := "0000000000000";	-- NOP
tmp(4) := "1001001000100";	-- JSR @SR_SET_LIMIT
tmp(5) := NOP & '0' & x"00"; 	 --%LABEL MAIN_LOOP
tmp(6) := "1001000101011";	-- JSR @SR_ATUALIZAR_DISPLAY
tmp(7) := "0000000000000";	-- NOP
tmp(8) := "1001011101111";	-- JSR @SR_VERIFICA_LIMITE
tmp(9) := "0000000000000";	-- NOP
tmp(10) := "1001010010010";	-- JSR @SR_INCREMENTO_CONTADOR
tmp(11) := "0000000000000";	-- NOP
tmp(12) := "0110000111110";	-- JMP @SR_VERIFICA_FPGA_RESET  	#-- Se for reset, volta pro loop inicial, caso contrario main loop
tmp(13) := "0000000000000";	-- NOP
tmp(14) := NOP & '0' & x"00"; 	 --%LABEL SR_INICIALIZACAO #-- ZERAR VALORES DA MEMORIA (INICIALIZACAO) - DANI
tmp(15) := "0100000000000";	-- LDI $0                               	# Carrega 0 no acumulador
tmp(16) := "0101000000000";	-- STA @ADDR_CTE0                       	# Seta a constate CTE0
tmp(17) := "0100000000001";	-- LDI $1                               	# Carrega 1 no acumulador 
tmp(18) := "0101000000001";	-- STA @ADDR_CTE1                       	# Seta a constante CTE1
tmp(19) := "0100000001001";	-- LDI $9                               	# Carrega 9 no acumulador 
tmp(20) := "0101000001001";	-- STA @ADDR_CTE9                       	# Seta a constante CTE9
tmp(21) := NOP & '0' & x"00"; 	 ---- Inicializar endereços de memória
tmp(22) := "0001000000000";	-- LDA @ADDR_CTE0                        	#-- Load cte 0
tmp(23) := "0101000001010";	-- STA @ADDR_COUNTER_UNIDADE        
tmp(24) := "0101000001011";	-- STA @ADDR_COUNTER_DEZENA         
tmp(25) := "0101000001100";	-- STA @ADDR_COUNTER_CENTENA        
tmp(26) := "0101000001101";	-- STA @ADDR_COUNTER_MILHAR         
tmp(27) := "0101000001110";	-- STA @ADDR_COUNTER_DEZ_MILHAR     
tmp(28) := "0101000001111";	-- STA @ADDR_COUNTER_CEN_MILHAR     
tmp(29) := "0101000010000";	-- STA @ADDR_LIMIT_COUNTER_UNIDADE  
tmp(30) := "0101000010001";	-- STA @ADDR_LIMIT_COUNTER_DEZENA   
tmp(31) := "0101000010010";	-- STA @ADDR_LIMIT_COUNTER_CENTENA  
tmp(32) := "0101000010011";	-- STA @ADDR_LIMIT_COUNTER_MILHAR   
tmp(33) := "0101000010100";	-- STA @ADDR_LIMIT_COUNTER_DEZ_MILHAR
tmp(34) := "0101000010101";	-- STA @ADDR_LIMIT_COUNTER_CEN_MILHAR
tmp(35) := "0101000010110";	-- STA @ADDR_FLAG_OVERFLOW
tmp(36) := "0101000010111";	-- STA @ADDR_FLAG_INIBICAO
tmp(37) := "0101101100100";	-- STA @FPGA_RESET
tmp(38) := "0101111111111";	-- STA @CLEAR_KEY0
tmp(39) := "0101111111110";	-- STA @CLEAR_KEY1
tmp(40) := "0101100000000";	-- STA @LEDR
tmp(41) := "1010000000000";	-- RET @ADDR_CTE0                      	#-- Exit inicialization sub routine
tmp(42) := "0000000000000";	-- NOP                                 	#-- === FIM INICIALIZAR CTE's  ===
tmp(43) := NOP & '0' & x"00"; 	 --%LABEL SR_ATUALIZAR_DISPLAY #-- ATUALIZAR DISPLAY - DANI
tmp(44) := "0001000001010";	-- LDA  @ADDR_COUNTER_UNIDADE    	#-- LOAD UNIDADE
tmp(45) := "0101100100000";	-- STA  @HEX0                    	#-- ARMAZENA EM HEX0
tmp(46) := "0001000001011";	-- LDA  @ADDR_COUNTER_DEZENA     	#-- LOAD DEZENA 
tmp(47) := "0101100100001";	-- STA  @HEX1                    	#-- ARMAZENA EM HEX1
tmp(48) := "0001000001100";	-- LDA  @ADDR_COUNTER_CENTENA    	#-- LOAD CENTENA
tmp(49) := "0101100100010";	-- STA  @HEX2                    	#-- ARMAZENA EM HEX2
tmp(50) := "0001000001101";	-- LDA  @ADDR_COUNTER_MILHAR     	#-- LOAD MILHAR
tmp(51) := "0101100100011";	-- STA  @HEX3                    	#-- ARMAZENA EM HEX3
tmp(52) := "0001000001110";	-- LDA  @ADDR_COUNTER_DEZ_MILHAR 	#-- LOAD DEZ.MILHAR 
tmp(53) := "0101100100100";	-- STA  @HEX4                    	#-- ARMAZENA EM HEX4
tmp(54) := "0001000001111";	-- LDA  @ADDR_COUNTER_CEN_MILHAR 	#-- LOAD CEN.MILHAR 
tmp(55) := "0101100100101";	-- STA  @HEX5                    	#-- ARMAZENA EM HEX5
tmp(56) := NOP & '0' & x"00"; 	 ---- ATUALIZA LEDS OVERFLOW, INIBICAO
tmp(57) := "0001000010110";	-- LDA @ADDR_FLAG_OVERFLOW       	#-- LOAD FLAG OVERFLOW
tmp(58) := "0101100000001";	-- STA @LED_F_OVERFLOW           	#-- ARMAZENA NO LED
tmp(59) := "0001000010111";	-- LDA @ADDR_FLAG_INIBICAO       	#-- LOAD FLAG INIBICAO
tmp(60) := "0101100000001";	-- STA @LED_F_OVERFLOW           	#-- ARMAZENA NO LED
tmp(61) := "1010000000000";	-- RET @0                        	#-- EXIT SUB ROUTINE;
tmp(62) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_FPGA_RESET
tmp(63) := "0001101100100";	-- LDA @FPGA_RESET
tmp(64) := "1000000000000";	-- CEQ @ADDR_CTE0
tmp(65) := "0111000000001";	-- JEQ @LOOP_INICIAL                     	#Se reset fpga == 0 (está invertido), recomeça tudo
tmp(66) := "0000000000000";	-- NOP
tmp(67) := "0110000000101";	-- JMP @MAIN_LOOP    
tmp(68) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT             #-- CONFIGURAR LIMITE CONTADOR
tmp(69) := "0001000000001";	-- LDA @ADDR_CTE1                  	# LOAD CTE1 (explicito)
tmp(70) := "0101100000000";	-- STA @LEDR                       	# Acender o primeiro LED
tmp(71) := "0001101000000";	-- LDA @SWR                        	# Carrega valores dos SW
tmp(72) := "0101000010000";	-- STA @ADDR_LIMIT_COUNTER_UNIDADE 	# SET UNIDADE LIMIT
tmp(73) := "0101100100000";	-- STA @HEX0                       	# Mostra o valor escolhido em HEX0
tmp(74) := "0001101100001";	-- LDA @KEY1                       	# LOAD KEY1
tmp(75) := "1000000000001";	-- CEQ @ADDR_CTE1                  	# KEY1 == 1
tmp(76) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(77) := "0111001010000";	-- JEQ @SR_SET_LIMIT_DEZ           	# If Key1 apertado: jmp configurar limite dezena
tmp(78) := "0000000000000";	-- NOP
tmp(79) := "0110001000100";	-- JMP @SR_SET_LIMIT           
tmp(80) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT_DEZ
tmp(81) := "0100000000010";	-- LDI $2                          	# LOAD 2 (explicito)
tmp(82) := "0101100000000";	-- STA @LEDR                       	# Acender o segundo LED
tmp(83) := "0001101000000";	-- LDA @SWR                        	# Carrega valores dos SW
tmp(84) := "0101000010001";	-- STA @ADDR_LIMIT_COUNTER_DEZENA  	# SET UNIDADE LIMIT
tmp(85) := "0101100100001";	-- STA @HEX1                       	# Mostra o valor escolhido em HEX1
tmp(86) := "0001101100001";	-- LDA @KEY1                       	# LOAD KEY1
tmp(87) := "1000000000001";	-- CEQ @ADDR_CTE1                  	# KEY1 == 1?
tmp(88) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(89) := "0111001011100";	-- JEQ @SR_SET_LIMIT_CENT          	# If Key1 apertado: jmp configurar limite CENT
tmp(90) := "0000000000000";	-- NOP
tmp(91) := "0110001010000";	-- JMP @SR_SET_LIMIT_DEZ           	# if key1 not apertado: refaz o processo para DEZENA
tmp(92) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT_CENT
tmp(93) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(94) := "0100000000100";	-- LDI $4                          	# LOAD 4 (explicito)
tmp(95) := "0101100000000";	-- STA @LEDR                       	# Acender o terceiro LED
tmp(96) := "0001101000000";	-- LDA @SWR                        	# Carrega valores dos SW
tmp(97) := "0101000010010";	-- STA @ADDR_LIMIT_COUNTER_CENTENA 	# SET CENTENA LIMIT
tmp(98) := "0101100100010";	-- STA @HEX2                       	# Mostra o valor escolhido em HEX2
tmp(99) := "0001101100001";	-- LDA @KEY1                       	# LOAD KEY1
tmp(100) := "1000000000001";	-- CEQ @ADDR_CTE1                  	# KEY1 == 1?
tmp(101) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(102) := "0111001101001";	-- JEQ @SR_SET_LIMIT_MILHAR        	# If Key1 apertado: jmp configurar limite MILHAR
tmp(103) := "0000000000000";	-- NOP
tmp(104) := "0110001011100";	-- JMP @SR_SET_LIMIT_CENT          	# if key1 not apertado: refaz o processo para CENTENA
tmp(105) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT_MILHAR
tmp(106) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(107) := "0100000001000";	-- LDI $8                          	# Load 8 (explicito)
tmp(108) := "0101100000000";	-- STA @LEDR                       	# Acender o 4 LED
tmp(109) := "0001101000000";	-- LDA @SWR                        	# Carrega valores dos SW
tmp(110) := "0101000010011";	-- STA @ADDR_LIMIT_COUNTER_MILHAR  	# SET UNIDADE LIMIT
tmp(111) := "0101100100011";	-- STA @HEX3                       	# Mostra o valor escolhido em HEX3
tmp(112) := "0001101100001";	-- LDA @KEY1                       	# LOAD KEY1
tmp(113) := "1000000000001";	-- CEQ @ADDR_CTE1                  	# KEY1 == 1?
tmp(114) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(115) := "0111001110110";	-- JEQ @SR_SET_LIMIT_DEZ_MILHAR    	# If Key1 apertado: jmp configurar limite DEZ_MILHAR
tmp(116) := "0000000000000";	-- NOP
tmp(117) := "0110001101001";	-- JMP @SR_SET_LIMIT_MILHAR        	# if key1 not apertado: refaz o processo para MILHAR
tmp(118) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT_DEZ_MILHAR
tmp(119) := "0101111111110";	-- STA @CLEAR_KEY1                    	# RESET KEY1
tmp(120) := "0100000010000";	-- LDI $16                            	# Load 16 (explicito)
tmp(121) := "0101100000000";	-- STA @LEDR
tmp(122) := "0001101000000";	-- LDA @SWR                           	# Carrega valores dos SW
tmp(123) := "0101000010100";	-- STA @ADDR_LIMIT_COUNTER_DEZ_MILHAR 	# SET DEZ_MILHAR LIMIT
tmp(124) := "0101100100100";	-- STA @HEX4                          	# Mostra o valor escolhido em HEX4
tmp(125) := "0001101100001";	-- LDA @KEY1                          	# LOAD KEY1
tmp(126) := "1000000000001";	-- CEQ @ADDR_CTE1                     	# KEY1 == 1?
tmp(127) := "0101111111110";	-- STA @CLEAR_KEY1                 	# RESET KEY1
tmp(128) := "0111010000011";	-- JEQ @SR_SET_LIMIT_CENT_MILHAR      	# If Key1 apertado: jmp configurar limite CENT_MILHAR
tmp(129) := "0000000000000";	-- NOP
tmp(130) := "0110001110110";	-- JMP @SR_SET_LIMIT_DEZ_MILHAR       	# if key1 not apertado: refaz o processo para MILHAR
tmp(131) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_LIMIT_CENT_MILHAR
tmp(132) := "0101111111110";	-- STA @CLEAR_KEY1                    	# RESET KEY1
tmp(133) := "0100000100000";	-- LDI $32                            	# Load 32 (explicito)
tmp(134) := "0101100000000";	-- STA @LEDR                          	# Acender o 6 LED
tmp(135) := "0001101000000";	-- LDA @SWR                           	# Carrega valores dos SW
tmp(136) := "0101000010101";	-- STA @ADDR_LIMIT_COUNTER_CEN_MILHAR 	# SET CENT_MILHAR LIMIT
tmp(137) := "0101100100101";	-- STA @HEX5                          	# Mostra o valor escolhido em HEX5
tmp(138) := "0001101100001";	-- LDA @KEY1                          	# LOAD KEY1
tmp(139) := "1000000000000";	-- CEQ @ADDR_CTE0                     	# KEY1 == 0? Se nao tiver clicado continua configurando, else terminou de configurar
tmp(140) := "0101111111110";	-- STA @CLEAR_KEY1                    	# RESET KEY1
tmp(141) := "0111010000011";	-- JEQ @SR_SET_LIMIT_CENT_MILHAR      	# If Key1 apertado: jmp configurar limite CENT_MILHAR
tmp(142) := "0000000000000";	-- NOP
tmp(143) := "0001000000000";	-- LDA @ADDR_CTE0                     
tmp(144) := "0101100000000";	-- STA @LEDR                          	# Reset LEDR, as the limit setting is completed
tmp(145) := "1010000000000";	-- RET $0
tmp(146) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_CONTADOR
tmp(147) := "0001101100000";	-- LDA  @KEY0                       	# Carrega KEY0
tmp(148) := "1000000000001";	-- CEQ  @ADDR_CTE1                  	# Key0 == 1?
tmp(149) := "0101111111111";	-- STA  @CLEAR_KEY0                 	# Reset key0
tmp(150) := "0111010011111";	-- JEQ  @SR_INCREMENTO_UNIDADE      	# If key0==1: incrementacontador
tmp(151) := "0000000000000";	-- NOP
tmp(152) := "1010000000000";	-- RET  $0
tmp(153) := "0001000010111";	-- LDA  @ADDR_FLAG_INIBICAO         	# LOAD FLAG INIBICAO
tmp(154) := "1000000000000";	-- CEQ  @ADDR_CTE0                  	# Inibicao == 0?
tmp(155) := "0111010011111";	-- JEQ  @SR_INCREMENTO_UNIDADE      	# IF inib == 0 : incrementa, else RET
tmp(156) := "0000000000000";	-- NOP
tmp(157) := "1010000000000";	-- RET  $0
tmp(158) := NOP & '0' & x"00"; 	 ---- 1) UNIDADE
tmp(159) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_UNIDADE
tmp(160) := "0001000001010";	-- LDA  @ADDR_COUNTER_UNIDADE 	#-- LOAD UNIDADE
tmp(161) := "1000000001001";	-- CEQ  @ADDR_CTE9            	#-- COMPARA COM 9
tmp(162) := "0111010101000";	-- JEQ  @SR_INCREMENTO_DEZENA 	#PULA PARA INCREMENTO DE DEZENA
tmp(163) := "0000000000000";	-- NOP
tmp(164) := NOP & '0' & x"00"; 	 ---- IF (UNIDADE != 9): {UNIDADE++} 
tmp(165) := "0010000000001";	-- SOMA @ADDR_CTE1            	#-- SOMA 1        
tmp(166) := "0101000001010";	-- STA  @ADDR_COUNTER_UNIDADE 	#-- SET UNIDADE += 1;
tmp(167) := "1010000000000";	-- RET  @ADDR_CTE0            	#-- EXIT SUB ROUTINE;
tmp(168) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_DEZENA
tmp(169) := NOP & '0' & x"00"; 	 ---- ELSE (UNIDADE == 9): {UNIDADE=0; DEZENA++}
tmp(170) := "0001000000000";	-- LDA  @ADDR_CTE0            	#-- LOAD CTE 0
tmp(171) := "0101000001010";	-- STA  @ADDR_COUNTER_UNIDADE 	#-- SET UNIDADE = 0 | RAM[10] - UNIDADE;
tmp(172) := NOP & '0' & x"00"; 	 ---- 2) DEZENA
tmp(173) := "0001000001011";	-- LDA  @ADDR_COUNTER_DEZENA  	#-- LOAD DEZENA 
tmp(174) := "1000000001001";	-- CEQ  @ADDR_CTE9            	#-- COMPARA COM 9
tmp(175) := "0111010110101";	-- JEQ  @SR_INCREMENTO_CENTENA 	#PULA PARA INCREMENTO DE CENTENA
tmp(176) := "0000000000000";	-- NOP
tmp(177) := NOP & '0' & x"00"; 	 ---- IF DEZENA != 9: {DEZENA++} 
tmp(178) := "0010000000001";	-- SOMA @ADDR_CTE1            	#-- SOMA 1       
tmp(179) := "0101000001011";	-- STA  @ADDR_COUNTER_DEZENA  	#-- SET DEZENA += 1;
tmp(180) := "1010000000000";	-- RET  @ADDR_CTE0            	#-- EXIT SUB ROUTINE;
tmp(181) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_CENTENA
tmp(182) := NOP & '0' & x"00"; 	 ---- ELSE (DEZENA == 9): {DEZENA=0; CENTENA++}
tmp(183) := "0001000000000";	-- LDA  @ADDR_CTE0            	#-- LOAD CTE 0
tmp(184) := "0101000001011";	-- STA  @ADDR_COUNTER_DEZENA  	#-- SET DEZENA = 0 
tmp(185) := NOP & '0' & x"00"; 	 ---- 3) CENTENA
tmp(186) := "0001000001100";	-- LDA  @ADDR_COUNTER_CENTENA  	#-- LOAD CENTENA 
tmp(187) := "1000000001001";	-- CEQ  @ADDR_CTE9             	#-- COMPARA COM 9 
tmp(188) := "0111011000010";	-- JEQ  @SR_INCREMENTO_MILHAR  	#PULA PARA INCREMENTO DE MILHAR
tmp(189) := "0000000000000";	-- NOP
tmp(190) := NOP & '0' & x"00"; 	 ---- IF CENTENA != 9: {CENTENA++} 
tmp(191) := "0010000000001";	-- SOMA @ADDR_CTE1             	#-- SOMA 1        
tmp(192) := "0101000001100";	-- STA  @ADDR_COUNTER_CENTENA  	#-- SET CENTENA += 1;
tmp(193) := "1010000000000";	-- RET  @ADDR_CTE0             	#-- EXIT SUB ROUTINE;
tmp(194) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_MILHAR -- ELSE (CENTENA == 9): {CENTENA=0; MILHAR++}
tmp(195) := "0001000000000";	-- LDA  @ADDR_CTE0             	#-- LOAD CTE 0
tmp(196) := "0101000001100";	-- STA  @ADDR_COUNTER_CENTENA  	#-- SET CENTENA = 0
tmp(197) := NOP & '0' & x"00"; 	 ---- 4) MILHARES
tmp(198) := "0001000001101";	-- LDA  @ADDR_COUNTER_MILHAR      	#-- LOAD MILHAR   
tmp(199) := "1000000001001";	-- CEQ  @ADDR_CTE9                	#-- COMPARA COM 9
tmp(200) := "0111011001110";	-- JEQ  @SR_INCREMENTO_DEZ_MILHAR 	#-- PULA PARA INCREMENTO DE DEZ MILHAR
tmp(201) := "0000000000000";	-- NOP
tmp(202) := NOP & '0' & x"00"; 	 ---- IF MILHAR != 9: {MILHAR++} 
tmp(203) := "0010000000001";	-- SOMA @ADDR_CTE1                	#-- SOMA 1        
tmp(204) := "0101000001101";	-- STA  @ADDR_COUNTER_MILHAR      	#-- SET MILHAR += 1;
tmp(205) := "1010000000000";	-- RET  @ADDR_CTE0                	#-- EXIT SUB ROUTINE;
tmp(206) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_DEZ_MILHAR -- ELSE (MILHAR == 9): {MILHAR=0; DEZ_MILHAR++}
tmp(207) := "0001000000000";	-- LDA  @ADDR_CTE0                	#-- LOAD CTE 0
tmp(208) := "0101000001101";	-- STA  @ADDR_COUNTER_MILHAR      	#-- SET MILHAR = 0 
tmp(209) := NOP & '0' & x"00"; 	 ---- 5) DEZ. MILHARES
tmp(210) := "0001000001110";	-- LDA  @ADDR_COUNTER_DEZ_MILHAR     	#-- LOAD DEZ.MILHAR   
tmp(211) := "1000000001001";	-- CEQ  @ADDR_CTE9                   	#-- COMPARA COM 9 
tmp(212) := "0111011011010";	-- JEQ  @SR_INCREMENTO_CEN_MILHAR    	#-- PULA PARA INCREMENTO DE CEN.MILHAR
tmp(213) := "0000000000000";	-- NOP
tmp(214) := NOP & '0' & x"00"; 	 ---- IF DEZ.MILHAR != 9: {DEZ.MILHAR++} 
tmp(215) := "0010000000001";	-- SOMA @ADDR_CTE1                   	#-- SOMA 1  
tmp(216) := "0101000001110";	-- STA  @ADDR_COUNTER_DEZ_MILHAR     	#-- SET DEZ.MILHAR += 1;
tmp(217) := "1010000000000";	-- RET  @ADDR_CTE0                   	#-- EXIT SUB ROUTINE;
tmp(218) := NOP & '0' & x"00"; 	 --%LABEL SR_INCREMENTO_CEN_MILHAR   #-- ELSE (DEZ.MILHAR == 9): {DEZ.MILHAR=0; CEN.MILHAR++}
tmp(219) := "0001000000000";	-- LDA  @ADDR_CTE0  	#-- LOAD CTE 0
tmp(220) := "0101000001110";	-- STA  @ADDR_COUNTER_DEZ_MILHAR     	#-- SET DEZ.MILHAR = 0 
tmp(221) := NOP & '0' & x"00"; 	 ---- 6) CEN. MILHARES
tmp(222) := "0001000001111";	-- LDA  @ADDR_COUNTER_CEN_MILHAR     	#-- LOAD CEN.MILHAR 
tmp(223) := "1000000001001";	-- CEQ  @ADDR_CTE9                   	#-- COMPARA COM 9 
tmp(224) := "0111011100111";	-- JEQ  @SR_SET_OVERFLOW 	#PULA PARA FLAG OVErFLOW E LIMITE ATINGIDO
tmp(225) := "0000000000000";	-- NOP
tmp(226) := NOP & '0' & x"00"; 	 ---- IF CEN.MILHAR != 9: {CEN.MILHAR++} 
tmp(227) := "0010000000001";	-- SOMA @ADDR_CTE1                   	#-- SOMA 1
tmp(228) := "0101000001111";	-- STA  @ADDR_COUNTER_CEN_MILHAR     	#-- SET CEN.MILHAR += 1;
tmp(229) := "1010000000000";	-- RET  @ADDR_CTE0                   	#-- EXIT SUB ROUTINE;
tmp(230) := NOP & '0' & x"00"; 	 ---- ELSE (CEN.MILHAR == 9): {CEN.MILHAR=10; OVERFLOW=1 INIBI=1}
tmp(231) := NOP & '0' & x"00"; 	 --%LABEL SR_SET_OVERFLOW         #-- OVERFLOW E INIBICAO
tmp(232) := "0001000001111";	-- LDA  @ADDR_COUNTER_CEN_MILHAR  	#-- LOAD CEN.MILHAR 
tmp(233) := "0010000000001";	-- SOMA @ADDR_CTE1                	#-- SOMA 1
tmp(234) := "0101000001111";	-- STA  @ADDR_COUNTER_CEN_MILHAR  	#-- SET CEN.MILHAR += 1;
tmp(235) := "0001000000001";	-- LDA  @ADDR_CTE1                	#-- LOAD CTE 1
tmp(236) := "0101000010111";	-- STA  @ADDR_FLAG_INIBICAO       	#-- FLAG_INIBICAO = 1
tmp(237) := "0101000010110";	-- STA  @ADDR_FLAG_OVERFLOW       	#-- FLAG_OVERFLOW = 1
tmp(238) := "1010000000000";	-- RET  @ADDR_CTE0                	#-- EXIT SUB ROUTINE - INCREMENTA;
tmp(239) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE -- SUB-ROTINA LIMITE: VERIFICAR SE ATINGIU O LIMITE - DANI
tmp(240) := NOP & '0' & x"00"; 	 ---- 1) CEN.MILHAR
tmp(241) := "0001000010101";	-- LDA @ADDR_LIMIT_COUNTER_CEN_MILHAR   	#-- LOAD LIMITE CEN.MILHAR
tmp(242) := "1000000001111";	-- CEQ @ADDR_COUNTER_CEN_MILHAR         	#-- VERIFY (COUNTER == LIMIT)
tmp(243) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(244) := "0111011110111";	-- JEQ @SR_VERIFICA_LIMITE_DEZ_MILHAR   	#-- Jump to next verification
tmp(245) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(246) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(247) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE_DEZ_MILHAR #-- 2) DEZ.MILHAR
tmp(248) := "0100000100000";	-- LDI $32 
tmp(249) := "0101100000000";	-- STA @LEDR                            	#-- Set LEDR[5] ON (limit_cent_milhar_atingido)
tmp(250) := "0001000010100";	-- LDA @ADDR_LIMIT_COUNTER_DEZ_MILHAR   	#-- LOAD LIMITE DEZ.MILHAR
tmp(251) := "1000000001110";	-- CEQ @ADDR_COUNTER_DEZ_MILHAR         	#-- VERIFY (COUNTER == LIMIT)
tmp(252) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(253) := "0111100000000";	-- JEQ @SR_VERIFICA_LIMITE_MILHAR       	#-- Jump to next verification
tmp(254) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(255) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(256) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE_MILHAR     #-- 3) MILHAR
tmp(257) := "0100000110000";	-- LDI $48
tmp(258) := "0101100000000";	-- STA @LEDR                            	# LEDR[5..4] ON - Limit cent_milhar and dez_milhar atingido
tmp(259) := "0001000010011";	-- LDA @ADDR_LIMIT_COUNTER_MILHAR       	#-- LOAD LIMITE MILHAR
tmp(260) := "1000000001101";	-- CEQ @ADDR_COUNTER_MILHAR             	#-- VERIFY (COUNTER == LIMIT)
tmp(261) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(262) := "0111100001001";	-- JEQ @SR_VERIFICA_LIMITE_CENTENA      	#-- Jump to next verification
tmp(263) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(264) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(265) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE_CENTENA    #-- 4) CENTENA
tmp(266) := "0100000111000";	-- LDI $56
tmp(267) := "0101100000000";	-- STA @LEDR                            	# LEDR[5..3] ON - Limit cent_milhar, dez_milhar, milhar atingido
tmp(268) := "0001000010010";	-- LDA @ADDR_LIMIT_COUNTER_CENTENA      	#-- LOAD LIMITE CENTENA
tmp(269) := "1000000001100";	-- CEQ @ADDR_COUNTER_CENTENA            	#-- VERIFY (COUNTER == LIMIT)
tmp(270) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(271) := "0111100010010";	-- JEQ @SR_VERIFICA_LIMITE_DEZENA       	#-- Jump to next verification
tmp(272) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(273) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(274) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE_DEZENA     #-- 5) DEZENA
tmp(275) := "0100000111100";	-- LDI $60
tmp(276) := "0101100000000";	-- STA @LEDR                            	# LEDR[5..2] ON - Limit cent_milhar, dez_milhar, milhar, cent atingido
tmp(277) := "0001000010001";	-- LDA @ADDR_LIMIT_COUNTER_DEZENA   	#-- LOAD LIMITE DEZENA
tmp(278) := "1000000001011";	-- CEQ @ADDR_COUNTER_DEZENA             	#-- VERIFY (COUNTER == LIMIT)
tmp(279) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(280) := "0111100011011";	-- JEQ @SR_VERIFICA_LIMITE_UNIDADE      	#-- Jump to next verification
tmp(281) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(282) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(283) := NOP & '0' & x"00"; 	 --%LABEL SR_VERIFICA_LIMITE_UNIDADE #-- 1) UNIDADE
tmp(284) := "0100000111110";	-- LDI $62
tmp(285) := "0101100000000";	-- STA @LEDR                            	# LEDR[5..1] ON - Limit cent_milhar, dez_milhar, milhar, cent, dez atingido
tmp(286) := "0001000010000";	-- LDA @ADDR_LIMIT_COUNTER_UNIDADE   	#-- LOAD LIMITE UNIDADE
tmp(287) := "1000000001010";	-- CEQ @ADDR_COUNTER_UNIDADE         	#-- VERIFY (COUNTER == LIMIT)
tmp(288) := NOP & '0' & x"00"; 	 ----  IF (COUNTER == LIMIT): {CONTINUE}
tmp(289) := "0111100100100";	-- JEQ @SR_ATINGIU_LIMITE            	#-- JUMP SR 'LIMITE ATINGIDO'
tmp(290) := NOP & '0' & x"00"; 	 ----  ELSE (COUNTER != LIMIT): {FLAG INIBICAO=FALSE}
tmp(291) := "0110100101010";	-- JMP @SR_NAO_ATINGIU_LIMITE           	#-- JUMP SR 'LIMITE NAO ATINGIDO'
tmp(292) := NOP & '0' & x"00"; 	 --%LABEL SR_ATINGIU_LIMITE             #-- SUB-ROTINA LIMITE A): MARCA LIMITE ATINGIDO - DANI
tmp(293) := "0001000000000";	-- LDA $0 
tmp(294) := "0101100000000";	-- STA @LEDR                            	#-- Clear LEDR, as limit has reached
tmp(295) := "0001000000001";	-- LDA @ADDR_CTE1                       	#-- LOAD CTE 1
tmp(296) := "0101000010111";	-- STA @ADDR_FLAG_INIBICAO              	#-- FLAG_INIBICAO = 1
tmp(297) := "1010000000000";	-- RET                                  	#-- EXIT COUNTER LIMIT VERIFICATION SUB-ROUTINE
tmp(298) := NOP & '0' & x"00"; 	 --%LABEL SR_NAO_ATINGIU_LIMITE         #-- SUB-ROTINA LIMITE B): MARCA LIMITE NÃO ATINGIDO - DANI
tmp(299) := "0001000000000";	-- LDA @ADDR_CTE0                       	#-- LOAD CTE 0
tmp(300) := "0101000010111";	-- STA @ADDR_FLAG_INIBICAO              	#-- FLAG_INIBICAO = 0
tmp(301) := "1010000000000";	-- RET                                  	#-- EXIT COUNTER LIMIT VERIFICATION SUB-ROUTINE

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;
