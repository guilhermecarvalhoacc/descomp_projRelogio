decoderbinario